`define PROGRAM "programs/add.mem"
`define MICROCODE "microcode.mem"
`define CONSTANTPOOL_ADDRESS 'h0048
`define LOCALVARIABLEFRAME_ADDRESS 'h0050
`define STACKPOINTER_ADDRESS 'h0060
