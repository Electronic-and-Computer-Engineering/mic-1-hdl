module uart_tb();

logic RX;
logic TX;

uart DUT(   .RX(RX),
            .TX(TX));
            
            
        
endmodule