module uart(
    input logic RX,
    
    output logic TX);
    

endmodule