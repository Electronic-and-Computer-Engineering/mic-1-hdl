`timescale 1 ns / 1 ps

module control_store (
    input [8:0] addr,
    input [