module tb_main_memory;

initial begin

end
endmodule 