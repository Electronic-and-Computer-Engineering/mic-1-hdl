`ifndef _mic1_include_
`define _mic1_include_

`define MIC1_PROGRAM "programs/add.mem"
`define MIC1_MICROCODE "microcode.mem"
`define CONSTANTPOOL_ADDRESS 'h0048
`define LOCALVARIABLEFRAME_ADDRESS 'h0050
`define STACKPOINTER_ADDRESS 'h0060
`define MEMORY_SIZE 'h0083

`endif
