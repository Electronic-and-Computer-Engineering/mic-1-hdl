module uart_rx(
    //INPUTS
    input logic clk,
    input logic baud,
    input logic rst,
    input logic data_in,
    //OUTPUTS
    output logic [7:0]data_out,
    output logic rx_done);
    

endmodule