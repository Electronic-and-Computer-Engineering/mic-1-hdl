module shifter( 
    // INPUTS
    input [31:0] ALU_out,
    input [1:0] Comand,
  
    // OUTPUTS
    output [31:0] Shifter_out,

   

endmodule