module decoder_tb(

    );
endmodule
