module tb_main-memory;

initial begin

end
endmodule 