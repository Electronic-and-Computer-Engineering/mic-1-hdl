`ifndef _mic1_include_
`define _mic1_include_

`define MIC1_PROGRAM "add.mem"
`define MIC1_MICROCODE "microcode.mem"
`define CONSTANTPOOL_ADDRESS 'h0048
`define LOCALVARIABLEFRAME_ADDRESS 'h004b
`define STACKPOINTER_ADDRESS 'h005b
`define MEMORY_SIZE 'h008b

`endif
