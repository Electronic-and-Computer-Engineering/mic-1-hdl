`timescale 1 ns / 1 ps

module mic1_tb;

initial begin
    $display("Hi");
    $finish;
end

endmodule
